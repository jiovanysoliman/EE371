
// Needs more work
module task2 (address, clock, data, wren, q);
logic [2:0] address [31:0];
logic input CLOCK_50;
logic input [9:0] SW;
logic output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;



endmodule 