// Top level module for lab 4
// Allows switching between task 1 and task 2 using SW[9]


module DE1_SoC(CLOCK_50, SW, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);


//// switch between task 1 and task 2. 
//Assign algo = SW[9];
//
//always_comb begin
//
//	case(SW[9]) begin
//	
//		0: counter counterAlgo ();
//	
//		1: binary binaryAlgo ();
//		
//	endcase
//
//
//end

//assign Start = ~KEY[3];
//assign Reset = ~KEY[0];

//seg7 LocOutMSB (.hex(Loc[4]), .leds(HEX1));
//seg7 LocOutLSB (.hex(Loc[3:0]), .leds(HEX0));

endmodule 