module binary #() (SW, Loc, Done, Found);

input logic [9:0] SW;
output logic [4:0] Loc;
output logic Done;
output logic Found;


endmodule 