module binary #(parameter InputWidth = 8, parameter LocWidth = 5) (CLOCK_50, A, Start, Reset, Loc, Done, Found);

input logic CLOCK_50;
input logic [InputWidth-1:0] A;
input logic Start;
input logic Reset;
output logic [LocWidth:0] Loc;
output logic Done;
output logic Found;





endmodule 	