module counter_toplevel();
endmodule 