module task2_toplevel ()

part1 task1 ();
part2 task2 ();

endmodule